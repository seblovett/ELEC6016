// cpu.sv
// Writen by seblovett
// Date Created Tue 18 Feb 2014 23:12:41 GMT
// <+Last Edited: Wed 26 Mar 2014 12:21:31 GMT by hl13g10 on hind.ecs.soton.ac.uk +>
//`include "options.sv"

module cpu #(parameter n = 8) ( //n - bus width
	input wire Clock, nReset, 
	input wire [9:0] SW,
`ifdef demo
	output logic [9:0] LED
`else
	output logic [7: 0] LED
`endif	
	);

timeunit 1ns; timeprecision 1ps;
import opcodes::*;

alu_functions_t AluOp;
PcSel_t PcSel;
logic[n-1:0] MemData;
wire [n-1:0] MemAddr; 
wire RegWe, WDataSel, AccStore, Op1Sel, ImmSel;

ram r (.Clock(Clock), .Address(MemAddr), .Data(MemData));

`ifdef demo
	always_comb
	begin
		case (opcodes_t'(MemData[7:4]))
			WAIT0: LED[9:8] = 2'b01;
			WAIT1: LED[9:8] = 2'b10;
			default: LED[9:8] = 2'b00;
		endcase
	end
`endif
control c 
(
	.Clock(Clock),
	.nReset(nReset),
	.RegWe(RegWe),
	.AluOp(AluOp),
	.OpCode(opcodes_t'(MemData[7:4])),
	.WDataSel(WDataSel),
	.PcSel(PcSel),
	.AccStore(AccStore),
	.Sw8(SW[8]),
	.Op1Sel(Op1Sel),
//	.Op2Sel(Op2Sel),
	.ImmSel(ImmSel)
);

datapath d
(
	.ImmSel(ImmSel),
	.MemData(MemData),
	.MemAddr(MemAddr),
	.Switches(SW[7:0]),
	.LEDs(LED[7:0]),
	.Clock(Clock),
	.nReset(nReset),
	.RegWe(RegWe),
	.AluOp(AluOp),
	.WDataSel(WDataSel),
	.PcSel(PcSel),
	.AccStore(AccStore),
	.Op1Sel(Op1Sel)
//	.Op2Sel(Op2Sel)
);


endmodule

