opcodes.sv