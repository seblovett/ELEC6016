//This is an options file to configure the processor

//demo adds some extra LED functionality to help.
//`define demo