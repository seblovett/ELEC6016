package opcodes;

// ALU funcitons

typedef enum logic [1:0] {ALU_ADD, ALU_MULT} alu_functions_t;

endpackage
